--****************************************************************
--Microsemi Corporation Proprietary and Confidential
--Copyright 2014 Microsemi Corporation.  All rights reserved
--
--ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
--ACCORDANCE WITH THE MICROSEMI LICENSE AGREEMENT AND MUST BE 
--APPROVED IN ADVANCE IN WRITING.
--
--Description: CoreCORDIC
--             CORDIC Word-serial Arctan LUT
--
--Rev:
--v4.0 12/2/2014  Porting in TGI framework
--
--SVN Revision Information:
--SVN$Revision:$
--SVN$Date:$
--
--Resolved SARS
--
--
--
--Notes:
--
--****************************************************************

-- This is an automatically generated file

-- CORDIC constant angle (arctan) LUT
LIBRARY IEEE;
  USE IEEE.std_logic_1164.all;
  USE IEEE.numeric_std.all;

ENTITY CORECORDIC_C0_CORECORDIC_C0_0_word_cROM IS
  GENERIC(
    LOGITER   : integer:=5;
    IN_BITS   : integer:=32;
    DP_BITS   : integer:=48  );
  PORT (iterCount : IN std_logic_vector(LOGITER-1 DOWNTO 0);
        arctan    : OUT std_logic_vector(DP_BITS-1 DOWNTO 0);
        rcprGain_fx : OUT std_logic_vector(IN_BITS-1 DOWNTO 0)  );
END ENTITY CORECORDIC_C0_CORECORDIC_C0_0_word_cROM;

ARCHITECTURE gen_rtl OF CORECORDIC_C0_CORECORDIC_C0_0_word_cROM IS
BEGIN
  PROCESS (iterCount)
  BEGIN
    CASE to_integer(unsigned(iterCount)) IS
      WHEN  0 => arctan <= "000100000000000000000000000000000000000000000000";
      WHEN  1 => arctan <= "000010010111001000000010100011101100111011111010";
      WHEN  2 => arctan <= "000001001111110110011100001011011010111101110010";
      WHEN  3 => arctan <= "000000101000100010001000111010100000111011101111";
      WHEN  4 => arctan <= "000000010100010110000110101000011000011100101100";
      WHEN  5 => arctan <= "000000001010001011101011111100001010110010000010";
      WHEN  6 => arctan <= "000000000101000101111011000011110010111000010100";
      WHEN  7 => arctan <= "000000000010100010111110001010101000100011101010";
      WHEN  8 => arctan <= "000000000001010001011111001010011010001101101000";
      WHEN  9 => arctan <= "000000000000101000101111100101110101110110011000";
      WHEN 10 => arctan <= "000000000000010100010111110011000000000001001001";
      WHEN 11 => arctan <= "000000000000001010001011111001100000101001010100";
      WHEN 12 => arctan <= "000000000000000101000101111100110000011001110000";
      WHEN 13 => arctan <= "000000000000000010100010111110011000001101100001";
      WHEN 14 => arctan <= "000000000000000001010001011111001100000110110101";
      WHEN 15 => arctan <= "000000000000000000101000101111100110000011011011";
      WHEN 16 => arctan <= "000000000000000000010100010111110011000001101110";
      WHEN 17 => arctan <= "000000000000000000001010001011111001100000110111";
      WHEN 18 => arctan <= "000000000000000000000101000101111100110000011011";
      WHEN 19 => arctan <= "000000000000000000000010100010111110011000001110";
      WHEN 20 => arctan <= "000000000000000000000001010001011111001100000111";
      WHEN 21 => arctan <= "000000000000000000000000101000101111100110000011";
      WHEN 22 => arctan <= "000000000000000000000000010100010111110011000010";
      WHEN 23 => arctan <= "000000000000000000000000001010001011111001100001";
      WHEN 24 => arctan <= "000000000000000000000000000101000101111100110000";
      WHEN 25 => arctan <= "000000000000000000000000000010100010111110011000";
      WHEN 26 => arctan <= "000000000000000000000000000001010001011111001100";
      WHEN 27 => arctan <= "000000000000000000000000000000101000101111100110";
      WHEN 28 => arctan <= "000000000000000000000000000000010100010111110011";
      WHEN 29 => arctan <= "000000000000000000000000000000001010001011111010";
      WHEN 30 => arctan <= "000000000000000000000000000000000101000101111101";
      WHEN 31 => arctan <= "000000000000000000000000000000000010100010111110";
      WHEN OTHERS => arctan <= (OTHERS=>'0');
    END CASE;
  END PROCESS;

  rcprGain_fx <= "00100110110111010011101101101010";

END ARCHITECTURE gen_rtl;

