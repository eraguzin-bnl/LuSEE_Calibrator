
-- This is an automatically generated file

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

package coreparameters IS
  constant ARCHITECT : integer := 1;
  constant MODE      : integer := 3;
  constant DP_OPTION : integer := 2;
  constant DP_WIDTH  : integer := 16;
  constant IN_BITS   : integer := 32;
  constant OUT_BITS  : integer := 32;
  constant ROUND     : integer := 3;
  constant COARSE    : integer := 1;
  constant ITERATIONS: integer := 32;
end coreparameters;
